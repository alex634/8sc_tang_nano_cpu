module instruction_rom
(
    input [7:0] addr,
    output reg [7:0] data
);

    always @ (addr) begin
        case (addr)
            0: data = 8'b11111111;
            1: data = 8'b11011111;
            2: data = 8'b11101111;
            3: data = 8'b11001110;
            4: data = 8'b10010010;
            5: data = 8'b10110000;
            6: data = 8'b11001101;
            7: data = 8'b10110000;
            8: data = 8'b11001100;
            9: data = 8'b10110000;
            10: data = 8'b11001011;
            11: data = 8'b10110000;
            12: data = 8'b11001010;
            13: data = 8'b10110000;
            14: data = 8'b11001001;
            15: data = 8'b10110000;
            16: data = 8'b11111111;
            17: data = 8'b11111111;
            18: data = 8'b11111111;
            19: data = 8'b11111111;
            20: data = 8'b11111111;
            21: data = 8'b11111111;
            22: data = 8'b11111111;
            23: data = 8'b11111111;
            24: data = 8'b11111111;
            25: data = 8'b11111111;
            26: data = 8'b11111111;
            27: data = 8'b11111111;
            28: data = 8'b11111111;
            29: data = 8'b11111111;
            30: data = 8'b11111111;
            31: data = 8'b11111111;
            32: data = 8'b11111111;
            33: data = 8'b11111111;
            34: data = 8'b11111111;
            35: data = 8'b11111111;
            36: data = 8'b11111111;
            37: data = 8'b11111111;
            38: data = 8'b11111111;
            39: data = 8'b11111111;
            40: data = 8'b11111111;
            41: data = 8'b11111111;
            42: data = 8'b11111111;
            43: data = 8'b11111111;
            44: data = 8'b11111111;
            45: data = 8'b11111111;
            46: data = 8'b11111111;
            47: data = 8'b11111111;
            48: data = 8'b11111111;
            49: data = 8'b11111111;
            50: data = 8'b11111111;
            51: data = 8'b11111111;
            52: data = 8'b11111111;
            53: data = 8'b11111111;
            54: data = 8'b11111111;
            55: data = 8'b11111111;
            56: data = 8'b11111111;
            57: data = 8'b11111111;
            58: data = 8'b11111111;
            59: data = 8'b11111111;
            60: data = 8'b11111111;
            61: data = 8'b11111111;
            62: data = 8'b11111111;
            63: data = 8'b11111111;
            64: data = 8'b11111111;
            65: data = 8'b11111111;
            66: data = 8'b11111111;
            67: data = 8'b11111111;
            68: data = 8'b11111111;
            69: data = 8'b11111111;
            70: data = 8'b11111111;
            71: data = 8'b11111111;
            72: data = 8'b11111111;
            73: data = 8'b11111111;
            74: data = 8'b11111111;
            75: data = 8'b11111111;
            76: data = 8'b11111111;
            77: data = 8'b11111111;
            78: data = 8'b11111111;
            79: data = 8'b11111111;
            80: data = 8'b11111111;
            81: data = 8'b11111111;
            82: data = 8'b11111111;
            83: data = 8'b11111111;
            84: data = 8'b11111111;
            85: data = 8'b11111111;
            86: data = 8'b11111111;
            87: data = 8'b11111111;
            88: data = 8'b11111111;
            89: data = 8'b11111111;
            90: data = 8'b11111111;
            91: data = 8'b11111111;
            92: data = 8'b11111111;
            93: data = 8'b11111111;
            94: data = 8'b11111111;
            95: data = 8'b11111111;
            96: data = 8'b11111111;
            97: data = 8'b11111111;
            98: data = 8'b11111111;
            99: data = 8'b11111111;
            100: data = 8'b11111111;
            101: data = 8'b11111111;
            102: data = 8'b11111111;
            103: data = 8'b11111111;
            104: data = 8'b11111111;
            105: data = 8'b11111111;
            106: data = 8'b11111111;
            107: data = 8'b11111111;
            108: data = 8'b11111111;
            109: data = 8'b11111111;
            110: data = 8'b11111111;
            111: data = 8'b11111111;
            112: data = 8'b11111111;
            113: data = 8'b11111111;
            114: data = 8'b11111111;
            115: data = 8'b11111111;
            116: data = 8'b11111111;
            117: data = 8'b11111111;
            118: data = 8'b11111111;
            119: data = 8'b11111111;
            120: data = 8'b11111111;
            121: data = 8'b11111111;
            122: data = 8'b11111111;
            123: data = 8'b11111111;
            124: data = 8'b11111111;
            125: data = 8'b11111111;
            126: data = 8'b11111111;
            127: data = 8'b11111111;
            128: data = 8'b11111111;
            129: data = 8'b11111111;
            130: data = 8'b11111111;
            131: data = 8'b11111111;
            132: data = 8'b11111111;
            133: data = 8'b11111111;
            134: data = 8'b11111111;
            135: data = 8'b11111111;
            136: data = 8'b11111111;
            137: data = 8'b11111111;
            138: data = 8'b11111111;
            139: data = 8'b11111111;
            140: data = 8'b11111111;
            141: data = 8'b11111111;
            142: data = 8'b11111111;
            143: data = 8'b11111111;
            144: data = 8'b11111111;
            145: data = 8'b11111111;
            146: data = 8'b11111111;
            147: data = 8'b11111111;
            148: data = 8'b11111111;
            149: data = 8'b11111111;
            150: data = 8'b11111111;
            151: data = 8'b11111111;
            152: data = 8'b11111111;
            153: data = 8'b11111111;
            154: data = 8'b11111111;
            155: data = 8'b11111111;
            156: data = 8'b11111111;
            157: data = 8'b11111111;
            158: data = 8'b11111111;
            159: data = 8'b11111111;
            160: data = 8'b11111111;
            161: data = 8'b11111111;
            162: data = 8'b11111111;
            163: data = 8'b11111111;
            164: data = 8'b11111111;
            165: data = 8'b11111111;
            166: data = 8'b11111111;
            167: data = 8'b11111111;
            168: data = 8'b11111111;
            169: data = 8'b11111111;
            170: data = 8'b11111111;
            171: data = 8'b11111111;
            172: data = 8'b11111111;
            173: data = 8'b11111111;
            174: data = 8'b11111111;
            175: data = 8'b11111111;
            176: data = 8'b11111111;
            177: data = 8'b11111111;
            178: data = 8'b11111111;
            179: data = 8'b11111111;
            180: data = 8'b11111111;
            181: data = 8'b11111111;
            182: data = 8'b11111111;
            183: data = 8'b11111111;
            184: data = 8'b11111111;
            185: data = 8'b11111111;
            186: data = 8'b11111111;
            187: data = 8'b11111111;
            188: data = 8'b11111111;
            189: data = 8'b11111111;
            190: data = 8'b11111111;
            191: data = 8'b11111111;
            192: data = 8'b11111111;
            193: data = 8'b11111111;
            194: data = 8'b11111111;
            195: data = 8'b11111111;
            196: data = 8'b11111111;
            197: data = 8'b11111111;
            198: data = 8'b11111111;
            199: data = 8'b11111111;
            200: data = 8'b11111111;
            201: data = 8'b11111111;
            202: data = 8'b11111111;
            203: data = 8'b11111111;
            204: data = 8'b11111111;
            205: data = 8'b11111111;
            206: data = 8'b11111111;
            207: data = 8'b11111111;
            208: data = 8'b11111111;
            209: data = 8'b11111111;
            210: data = 8'b11111111;
            211: data = 8'b11111111;
            212: data = 8'b11111111;
            213: data = 8'b11111111;
            214: data = 8'b11111111;
            215: data = 8'b11111111;
            216: data = 8'b11111111;
            217: data = 8'b11111111;
            218: data = 8'b11111111;
            219: data = 8'b11111111;
            220: data = 8'b11111111;
            221: data = 8'b11111111;
            222: data = 8'b11111111;
            223: data = 8'b11111111;
            224: data = 8'b11111111;
            225: data = 8'b11111111;
            226: data = 8'b11111111;
            227: data = 8'b11111111;
            228: data = 8'b11111111;
            229: data = 8'b11111111;
            230: data = 8'b11111111;
            231: data = 8'b11111111;
            232: data = 8'b11111111;
            233: data = 8'b11111111;
            234: data = 8'b11111111;
            235: data = 8'b11111111;
            236: data = 8'b11111111;
            237: data = 8'b11111111;
            238: data = 8'b11111111;
            239: data = 8'b11111111;
            240: data = 8'b11111111;
            241: data = 8'b11111111;
            242: data = 8'b11111111;
            243: data = 8'b11111111;
            244: data = 8'b11111111;
            245: data = 8'b11111111;
            246: data = 8'b11111111;
            247: data = 8'b11111111;
            248: data = 8'b11111111;
            249: data = 8'b11111111;
            250: data = 8'b11111111;
            251: data = 8'b11111111;
            252: data = 8'b11111111;
            253: data = 8'b11111111;
            254: data = 8'b11111111;
            255: data = 8'b11111111;
              
        endcase
    end

endmodule
